//// megafunction wizard: %RAM: 2-PORT%VBB%
//// GENERATION: STANDARD
//// VERSION: WM1.0
//// MODULE: altsyncram 
//
//// ============================================================
//// File Name: ram32x3port2.v
//// Megafunction Name(s):
//// 			altsyncram
////
//// Simulation Library Files(s):
//// 			altera_mf
//// ============================================================
//// ************************************************************
//// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
////
//// 17.0.0 Build 595 04/25/2017 SJ Lite Edition
//// ************************************************************
//
////Copyright (C) 2017  Intel Corporation. All rights reserved.
////Your use of Intel Corporation's design tools, logic functions 
////and other software and tools, and its AMPP partner logic 
////functions, and any output files from any of the foregoing 
////(including device programming or simulation files), and any 
////associated documentation or information are expressly subject 
////to the terms and conditions of the Intel Program License 
////Subscription Agreement, the Intel Quartus Prime License Agreement,
////the Intel MegaCore Function License Agreement, or other 
////applicable license agreement, including, without limitation, 
////that your use is for the sole purpose of programming logic 
////devices manufactured by Intel and sold by Intel or its 
////authorized distributors.  Please refer to the applicable 
////agreement for further details.
//
//module ram32x3port2 (
//	clock,
//	data,
//	rdaddress,
//	wraddress,
//	wren,
//	q);
//
//	input	  clock;
//	input	[2:0]  data;
//	input	[4:0]  rdaddress;
//	input	[4:0]  wraddress;
//	input	  wren;
//	output	[2:0]  q;
//`ifndef ALTERA_RESERVED_QIS
//// synopsys translate_off
//`endif
//	tri1	  clock;
//	tri0	  wren;
//`ifndef ALTERA_RESERVED_QIS
//// synopsys translate_on
//`endif
//
//endmodule
//
//// ============================================================
//// CNX file retrieval info
//// ============================================================
//// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
//// Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
//// Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
//// Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
//// Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
//// Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
//// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
//// Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
//// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
//// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "0"
//// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
//// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_B NUMERIC "0"
//// Retrieval info: PRIVATE: CLRdata NUMERIC "0"
//// Retrieval info: PRIVATE: CLRq NUMERIC "0"
//// Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
//// Retrieval info: PRIVATE: CLRrren NUMERIC "0"
//// Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
//// Retrieval info: PRIVATE: CLRwren NUMERIC "0"
//// Retrieval info: PRIVATE: Clock NUMERIC "0"
//// Retrieval info: PRIVATE: Clock_A NUMERIC "0"
//// Retrieval info: PRIVATE: Clock_B NUMERIC "0"
//// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
//// Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
//// Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "0"
//// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_B"
//// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
//// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
//// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
//// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
//// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
//// Retrieval info: PRIVATE: MEMSIZE NUMERIC "96"
//// Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "0"
//// Retrieval info: PRIVATE: MIFfilename STRING "ram32x3.mif"
//// Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "2"
//// Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
//// Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "1"
//// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "2"
//// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "2"
//// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
//// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "3"
//// Retrieval info: PRIVATE: REGdata NUMERIC "1"
//// Retrieval info: PRIVATE: REGq NUMERIC "1"
//// Retrieval info: PRIVATE: REGrdaddress NUMERIC "1"
//// Retrieval info: PRIVATE: REGrren NUMERIC "1"
//// Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
//// Retrieval info: PRIVATE: REGwren NUMERIC "1"
//// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
//// Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
//// Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
//// Retrieval info: PRIVATE: VarWidth NUMERIC "0"
//// Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "3"
//// Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "3"
//// Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "3"
//// Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "3"
//// Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
//// Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "0"
//// Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
//// Retrieval info: PRIVATE: enable NUMERIC "0"
//// Retrieval info: PRIVATE: rden NUMERIC "0"
//// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
//// Retrieval info: CONSTANT: ADDRESS_ACLR_B STRING "NONE"
//// Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK0"
//// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
//// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "BYPASS"
//// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_B STRING "BYPASS"
//// Retrieval info: CONSTANT: INIT_FILE STRING "ram32x3.mif"
//// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
//// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
//// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "32"
//// Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "32"
//// Retrieval info: CONSTANT: OPERATION_MODE STRING "DUAL_PORT"
//// Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
//// Retrieval info: CONSTANT: OUTDATA_REG_B STRING "CLOCK0"
//// Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
//// Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "M10K"
//// Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_MIXED_PORTS STRING "DONT_CARE"
//// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "5"
//// Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "5"
//// Retrieval info: CONSTANT: WIDTH_A NUMERIC "3"
//// Retrieval info: CONSTANT: WIDTH_B NUMERIC "3"
//// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
//// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
//// Retrieval info: USED_PORT: data 0 0 3 0 INPUT NODEFVAL "data[2..0]"
//// Retrieval info: USED_PORT: q 0 0 3 0 OUTPUT NODEFVAL "q[2..0]"
//// Retrieval info: USED_PORT: rdaddress 0 0 5 0 INPUT NODEFVAL "rdaddress[4..0]"
//// Retrieval info: USED_PORT: wraddress 0 0 5 0 INPUT NODEFVAL "wraddress[4..0]"
//// Retrieval info: USED_PORT: wren 0 0 0 0 INPUT GND "wren"
//// Retrieval info: CONNECT: @address_a 0 0 5 0 wraddress 0 0 5 0
//// Retrieval info: CONNECT: @address_b 0 0 5 0 rdaddress 0 0 5 0
//// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
//// Retrieval info: CONNECT: @data_a 0 0 3 0 data 0 0 3 0
//// Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
//// Retrieval info: CONNECT: q 0 0 3 0 @q_b 0 0 3 0
//// Retrieval info: GEN_FILE: TYPE_NORMAL ram32x3port2.v TRUE
//// Retrieval info: GEN_FILE: TYPE_NORMAL ram32x3port2.inc FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL ram32x3port2.cmp FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL ram32x3port2.bsf FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL ram32x3port2_inst.v FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL ram32x3port2_bb.v TRUE
//// Retrieval info: LIB_FILE: altera_mf
