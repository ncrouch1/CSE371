module FIFO_filter #(Size=10)();

endmodule
